library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


entity lutsIntelDP is
  Port ( 
    a2 : in unsigned(2 downto 0);
	b : in unsigned(5 downto 0);
	a2b0 : out unsigned(7 downto 0);
	b2 : out unsigned(5 downto 0));
end lutsIntelDP;


architecture rtl of lutsIntelDP is

signal combi : unsigned(5 downto 0);

begin

combi <= a2 & b(5 downto 3); 


with combi select a2b0 <=
"00000000" when "000000", 
"00000000" when "000001", 
"00000000" when "000010", 
"00000000" when "000011", 
"00000000" when "000100", 
"00000000" when "000101", 
"00000000" when "000110", 
"00000000" when "000111", 
"00000000" when "001000", 
"00000011" when "001001", 
"00000110" when "001010", 
"00001001" when "001011", 
"00001100" when "001100", 
"00001111" when "001101", 
"00010010" when "001110", 
"00010101" when "001111", 
"00000000" when "010000", 
"00000110" when "010001", 
"00001100" when "010010", 
"00010010" when "010011", 
"00011000" when "010100", 
"00011110" when "010101", 
"00100100" when "010110", 
"00101010" when "010111", 
"00000000" when "011000", 
"00001001" when "011001", 
"00010010" when "011010", 
"00011011" when "011011", 
"00100100" when "011100", 
"00101101" when "011101", 
"00110110" when "011110", 
"00111111" when "011111", 
"00000000" when "100000", 
"00001100" when "100001", 
"00011000" when "100010", 
"00100100" when "100011", 
"00110000" when "100100", 
"00111100" when "100101", 
"01001000" when "100110", 
"01010100" when "100111", 
"00000000" when "101000", 
"00001111" when "101001", 
"00011110" when "101010", 
"00101101" when "101011", 
"00111100" when "101100", 
"01001011" when "101101", 
"01011010" when "101110", 
"01101001" when "101111", 
"00000000" when "110000", 
"00010010" when "110001", 
"00100100" when "110010", 
"00110110" when "110011", 
"01001000" when "110100", 
"01011010" when "110101", 
"01101100" when "110110", 
"01111110" when "110111", 
"00000000" when "111000", 
"00010101" when "111001", 
"00101010" when "111010", 
"00111111" when "111011", 
"01010100" when "111100", 
"01101001" when "111101", 
"01111110" when "111110", 
"10010011" when others; 


with b select b2 <=
"000000" when "000000", 
"000000" when "000001", 
"000000" when "000010", 
"000000" when "000011", 
"000000" when "000100", 
"000000" when "000101", 
"000000" when "000110", 
"000000" when "000111", 
"000001" when "001000", 
"000001" when "001001", 
"000001" when "001010", 
"000001" when "001011", 
"000010" when "001100", 
"000010" when "001101", 
"000011" when "001110", 
"000011" when "001111", 
"000100" when "010000", 
"000100" when "010001", 
"000101" when "010010", 
"000101" when "010011", 
"000110" when "010100", 
"000110" when "010101", 
"000111" when "010110", 
"001000" when "010111", 
"001001" when "011000", 
"001001" when "011001", 
"001010" when "011010", 
"001011" when "011011", 
"001100" when "011100", 
"001101" when "011101", 
"001110" when "011110", 
"001111" when "011111", 
"010000" when "100000", 
"010001" when "100001", 
"010010" when "100010", 
"010011" when "100011", 
"010100" when "100100", 
"010101" when "100101", 
"010110" when "100110", 
"010111" when "100111", 
"011001" when "101000", 
"011010" when "101001", 
"011011" when "101010", 
"011100" when "101011", 
"011110" when "101100", 
"011111" when "101101", 
"100001" when "101110", 
"100010" when "101111", 
"100100" when "110000", 
"100101" when "110001", 
"100111" when "110010", 
"101000" when "110011", 
"101010" when "110100", 
"101011" when "110101", 
"101101" when "110110", 
"101111" when "110111", 
"110001" when "111000", 
"110010" when "111001", 
"110100" when "111010", 
"110110" when "111011", 
"111000" when "111100", 
"111010" when "111101", 
"111100" when "111110", 
"111110" when others;  


end rtl;
